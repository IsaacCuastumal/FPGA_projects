library verilog;
use verilog.vl_types.all;
entity easy_verilog_example is
end easy_verilog_example;
