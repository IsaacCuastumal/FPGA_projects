library verilog;
use verilog.vl_types.all;
entity testbench_4bit_adder is
end testbench_4bit_adder;
