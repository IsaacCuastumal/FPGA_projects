library verilog;
use verilog.vl_types.all;
entity tb_decoder_4to16 is
end tb_decoder_4to16;
