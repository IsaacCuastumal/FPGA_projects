library verilog;
use verilog.vl_types.all;
entity easy_vector_example is
end easy_vector_example;
