library verilog;
use verilog.vl_types.all;
entity literal_values is
end literal_values;
