library verilog;
use verilog.vl_types.all;
entity tb_shift_reg_pipo is
end tb_shift_reg_pipo;
