library verilog;
use verilog.vl_types.all;
entity tb_shift_reg_siso is
end tb_shift_reg_siso;
