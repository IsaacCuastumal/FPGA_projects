library verilog;
use verilog.vl_types.all;
entity waveforms is
end waveforms;
