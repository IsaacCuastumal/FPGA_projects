library verilog;
use verilog.vl_types.all;
entity tb_hex_7seg_decoder is
end tb_hex_7seg_decoder;
