module hello_world();

initial begin
 $display("\n\t My name is Isaac and I start the course today 05/FEB/2025! \n");
 
 end
 
 endmodule 