library verilog;
use verilog.vl_types.all;
entity bitwise_operators is
end bitwise_operators;
