library verilog;
use verilog.vl_types.all;
entity procedures is
end procedures;
