library verilog;
use verilog.vl_types.all;
entity my_first_testbench is
end my_first_testbench;
